
`ifndef RST_UVC_PKG_SV
`define RST_UVC_PKG_SV

`include "rst_uvc_if.sv"

package rst_uvc_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "rst_uvc_common.sv"
`include "rst_uvc_agent_cfg.sv"
`include "rst_uvc_cfg.sv"
`include "rst_uvc_item.sv"
`include "rst_uvc_driver.sv"
`include "rst_uvc_sequencer.sv"
`include "rst_uvc_monitor.sv"
`include "rst_uvc_cov.sv"
`include "rst_uvc_agent.sv"
`include "rst_uvc_env.sv"
`include "rst_uvc_sequence_lib.sv"

endpackage : rst_uvc_pkg

`endif // RST_UVC_PKG_SV
